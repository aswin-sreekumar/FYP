// Register file block

module Register_File(clk,rst,WE3,WD3,A1,A2,A3,RD1,RD2);

    input clk,rst,WE3;
    input [4:0]A1,A2,A3;
    input [31:0]WD3;
    output [31:0]RD1,RD2;

    reg [31:0] Register [31:0];

    always @ (posedge clk)
    begin
        if(WE3)
            Register[A3] <= WD3;
    end

    assign RD1 = (~rst) ? 32'd0 : Register[A1];
    assign RD2 = (~rst) ? 32'd0 : Register[A2];

    initial begin
        Register[0] = 32'h00000005;
        Register[1] = 32'h00000003;
        Register[2] = 32'h00000100;
        
        $monitor("\ntime = %d\n", $time, 
        "\tRegister[0] = %b\n", Register[0],   
        "\tRegister[1] = %b\n", Register[1],
        "\tRegister[2] = %b\n", Register[2]);

    end

endmodule