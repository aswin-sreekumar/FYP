// Recovery unit module

module Recovery_Unit(
    
);

endmodule