// MUX for ALU input and data memory to register
// Instantiated twice in top level

module Mux (a,b,s,c);

    input [31:0]a,b;
    input s;
    output [31:0]c;

    assign c = (~s) ? a : b ;
    
endmodule